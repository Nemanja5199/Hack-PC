module I_Gate(output[15:0] Y, input[15:0] A,B);
  

  
 assign Y= A&B;
  
 
endmodule 