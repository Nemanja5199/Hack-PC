

module ASCIItoData(output[15:0] A, input [7:0]B);




assign A = {8'b00000000,B};



endmodule